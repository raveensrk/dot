    function void print;
        $display("i_e = %p", i_e);
    endfunction: print
