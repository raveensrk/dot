function void build_phase(uvm_phase phase);
	super.build_phase(phase);
endfunction
