`uvm_fatal(get_name(), $sformatf("var = %0d", var));
