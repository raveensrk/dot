uvm_config_db#(int)::set(null, "db_name", "var_name", 1/*set value*/);
