if (expression) begin
end else begin
end
