fd = $fopen("file.log", "w");
