$fdisplay(fd, "%m: %s", "String");
