foreach (array[index]) begin
    $display("%s = %0d", index, array[index]);
end
