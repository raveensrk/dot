uvm_config_db#(int)::get(null, "db_name", "var_name", get_value);
