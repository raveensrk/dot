`ifdef DEBUG
`endif
