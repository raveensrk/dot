`uvm_error(get_name(), $sformatf("var = %0d", var));
