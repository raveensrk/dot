for (int i=0; i<=n; i++) begin
end
