case(sel)
    default: out = 0;
    2'b00: out = a;
    2'b01: out = b;
    2'b10: out = c;
endcase
